`timescale 1ns/1ps

module INSTRUCTION_FETCH(
	clk,
	rst,
	jump,
	branch,
	jump_addr,
	branch_addr,

	PC,
	IR
);

input clk, rst, jump, branch;
input [31:0] jump_addr, branch_addr;

output reg 	[31:0] PC;
output reg 	[31:0] IR;

reg [31:0] instruction [0:127];	// 127:0

// Instruction DM initialilation	// initial to always -> reset function
always @ (posedge clk or posedge rst) begin	
	if(rst) begin
	/*=================================================     連加     =================================================*/
		//$0 = 0, $1 = 1, $2 = 2, $3 = 3, $4 = 5, $5 = input, ($6,$7) = limit, $8 = TF, ($9,$10) = approx, ($25,$26) = ans
		instruction[ 0] = 32'b100011_00000_00101_00000_00000_000000;	// lw $5, 0($0)
		instruction[ 1] = 32'b000000_00000_00011_00110_00000_100000;	// add $6, $0, $3   
		instruction[ 2] = 32'b000000_00000_00011_00111_00000_100000;	// add $7, $0, $3        
		instruction[ 3] = 32'b101011_00000_00010_00000_00000_000001;	// sw $2, 1($0)		tmp answer: 2 
		instruction[ 4] = 32'b000000_00101_00001_01001_00000_100100;	// and $9, $5, $1   even or odd	  pc: 10
		instruction[ 5] = 32'b000101_00101_00011_00000_00000_000111;	// bne $5, $3, 7	special case: 3	(loop) 
		/*	Input == 3	*/
		instruction[ 6] = 32'b101011_00000_00100_00000_00000_000010;	// sw $4, 2($0)		tmp answer: 5
		instruction[ 7] = 32'b000000_00000_00000_00000_00000_100000;	// NOP 
		instruction[ 8] = 32'b000000_00001_01001_01001_00000_100010;	// sub $9, $1, $9                   20
		instruction[ 9] = 32'b000010_00000_00000_00000_00001_111011; 	// j  exit (123)                 
		instruction[10] = 32'b000000_00000_00000_00000_00000_100000;	// NOP                          
		instruction[11] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                           
		instruction[12] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                 30
		/*	loop (calculate n^-2)	*/
		instruction[13] = 32'b000000_00110_00101_01000_00000_101010;	// slt $8, $6, $5
		instruction[14] = 32'b000000_00000_00000_00000_00000_100000;	// NOP		                        
		instruction[15] = 32'b000000_00000_00000_00000_00000_100000;	// NOP                          
		instruction[16] = 32'b000000_00110_00111_00110_00000_100000; 	// add $6, $6, $7   				  40          
		instruction[17] = 32'b000100_01000_00000_00000_00000_001000; 	// beq $8, $0, 8                
		instruction[18] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                         
		instruction[19] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                       
		instruction[20] = 32'b000000_00110_00111_00110_00000_100000; 	// add $6, $6, $7                     50
		instruction[21] = 32'b000000_00111_00001_00111_00000_100000; 	// add $7, $7, $1               
		instruction[22] = 32'b000010_00000_00000_00000_00000_001101; 	// j 13	(loop)                   
		instruction[23] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                          
		instruction[24] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                60                     
		instruction[25] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                           
		/*	A($25) < x, B($26) > x	*/
		instruction[26] = 32'b000000_00101_01001_11001_00000_100000; 	// add $25, $5, $9  X<A                         
		instruction[27] = 32'b000000_00101_01001_11010_00000_100010; 	// sub $26, $5, $9  X>A
		instruction[28] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                70                           
		/*	cmpA	*/
		instruction[29] = 32'b000000_00000_00011_01001_00000_100000; 	// add $9, $0, $3
		instruction[30] = 32'b000000_11001_00010_11001_00000_100010; 	// sub $25, $25, $2
		instruction[31] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[32] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                80
		/*	cmpA1	*/
		instruction[33] = 32'b000000_01001_00111_01000_00000_101010; 	// slt $8, $9, $7   			      84
		instruction[34] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[35] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[36] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                90
		instruction[37] = 32'b000100_01000_00000_00000_00000_100101; 	// beq $8, $0, 37	(ansA)
		instruction[38] = 32'b000000_01001_01001_00110_00000_100000; 	// add $6, $9, $9
		instruction[39] = 32'b000000_11001_00000_01010_00000_100000; 	// add $10, $25, $0
		instruction[40] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                A0
 		instruction[41] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[42] = 32'b000000_00110_00110_00110_00000_100000; 	// add $6, $6, $6
		instruction[43] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
 		instruction[44] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                B0
		instruction[45] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		/*	cmpA2	*/
		instruction[46] = 32'b000000_01010_00110_01010_00000_100010; 	// sub $10, $10, $6
		instruction[47] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[48] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                C0
		instruction[49] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[50] = 32'b000000_01001_01010_01000_00000_101010; 	// slt $8, $9, $10
		instruction[51] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[52] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                D0
		instruction[53] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[54] = 32'b000101_01000_00000_11111_11111_110111; 	// bne $8, $0, -9	(cmp2)
		instruction[55] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[56] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                E0
		instruction[57] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[58] = 32'b000100_01010_01001_11111_11111_100010;	// beq $10, $9, -30	(cmp)
		instruction[59] = 32'b000000_01001_01010_01010_00000_100000; 	// add $10, $10, $9
		instruction[60] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                F0
		instruction[61] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[62] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[63] = 32'b000100_01010_00000_11111_11111_011101; 	// beq $10, $0, -35	(cmp)
		instruction[64] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                100
		instruction[65] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                            
		instruction[66] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[67] = 32'b000000_01001_00010_01001_00000_100000; 	// add $9, $9, $2
		instruction[68] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                110
		instruction[69] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[70] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[71] = 32'b000010_00000_00000_00000_00000_100001; 	// j 33	(comp1)
		instruction[72] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                120
		instruction[73] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[74] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		/*	ansA	*/
		instruction[75] = 32'b101011_00000_11001_00000_00000_000001; 	// sw $25, 1($0)
		/*	compB	*/
		instruction[76] = 32'b000000_00000_00011_01001_00000_100000; 	// add $9, $0, $3                     130
		instruction[77] = 32'b000000_11010_00010_11010_00000_100000; 	// add $26, $26, $2
		instruction[78] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[79] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                 
		/*	comp1B	*/               
		instruction[80] = 32'b000000_01001_00111_01000_00000_101010; 	// slt $8, $9, $7          			  140
		instruction[81] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[82] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[83] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[84] = 32'b000100_01000_00000_00000_00000_100101; 	// beq $8, $0, 37   (ansB)            150
		instruction[85] = 32'b000000_01001_01001_00110_00000_100000; 	// add $6, $9, $9
		instruction[86] = 32'b000000_11010_00000_01010_00000_100000; 	// add $10, $26, $0
		instruction[87] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                160
 		instruction[88] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[89] = 32'b000000_00110_00110_00110_00000_100000; 	// add $6, $6, $6 
		instruction[90] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
 		instruction[91] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[92] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		/*	comp2B	*/
		instruction[93] = 32'b000000_01010_00110_01010_00000_100010; 	// sub $10, $10, $6
		instruction[94] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[95] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[96] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[97] = 32'b000000_01001_01010_01000_00000_101010; 	// slt $8, $9, $10
		instruction[98] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[99] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[100] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[101] = 32'b000101_01000_00000_11111_11111_110111; 	// bne $8, $0, -9	(comp2B)
		instruction[102] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[103] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[104] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[105] = 32'b000100_01010_01001_11111_11111_100010; 	// beq $10, $9, -30	(compB)
		instruction[106] = 32'b000000_01010_01001_01010_00000_100000; 	// add $10, $10, $9
		instruction[107] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[108] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[109] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[110] = 32'b000100_01010_00000_11111_11111_011101; 	// beq $10, $0, -35 (compB)
		instruction[111] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[112] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                            
		instruction[113] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[114] = 32'b000000_01001_00010_01001_00000_100000; 	// add $9, $9, $2
		instruction[115] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[116] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[117] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		instruction[118] = 32'b000010_00000_00000_00000_00001_010000; 	// j 80	(comp1B)
		instruction[119] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[120] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[121] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP
		/*	ansB	*/
		instruction[122] = 32'b101011_00000_11010_00000_00000_000010; 	// sw $26, 2($0)
		instruction[123] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[124] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP                                
		instruction[125] = 32'b000000_00000_00000_00000_00000_100000; 	// NOP

		//for (i=126; i<128; i=i+1)  instruction[ i] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	end
	else begin
		if (PC[10:2] <= 8'd125)
			IR <= instruction[PC[10:2]]; //(0, 4, 8, ...) => (0, 1, 2, ...)
	end
end

// output program counter
always @(posedge clk or posedge rst)
begin
	if(rst)
		PC <= 32'd0;
	else begin
		if(PC[10:2] < 8'd125)
			PC <= (branch) ? branch_addr : ( (jump) ? jump_addr : (PC+4));
	end
end

endmodule